`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/07/2025 11:24:39 AM
// Design Name: 
// Module Name: twobitcounter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module twobitcounter(
    input clk, 
    output [1:0] Q
    );
    reg [1:0] temp=0;
    always @(posedge clk)
    begin
        temp = temp + 1;
    end
    assign Q = temp;
    
    
endmodule
